module top();

endmodule
module tb;

endmodule